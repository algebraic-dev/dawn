module registers(clock, read1, read2, data1, data2, reg_write, wrreg, wrdata);
    input wire clock;
endmodule